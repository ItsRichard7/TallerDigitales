module StateMachine ()

endmodule