module StateMachine (
	output logic rst, clk
);

Clock clock(
	.clk(clk)
);

endmodule