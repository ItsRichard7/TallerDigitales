module decoder (input v,x,y,z output a,b,c,d,e,f,g)

endmodule