module Battleship ()

endmodule