module Battleship_tb ()


endmodule