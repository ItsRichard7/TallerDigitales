module Clock_tb;

logic clk;

Clock clock(
	.clk(clk)
	);

endmodule